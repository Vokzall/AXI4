`ifndef AXI_DEFINES
`define AXI_DEFINES

`define AXI_ADDR_WIDTH 32
`define AXI_DATA_WIDTH 32
`define AXI_ID_WIDTH   4
`define AXI_STRB_WIDTH (`AXI_DATA_WIDTH/8)

`endif